`include "dat.vh"

module addattest;

	addat addat0(adclk, adsfl, advs, adhs, adfield, addat, inde, indat);

endmodule
